library ieee;
use ieee.std_logic_1164.all;

entity ff_d_14 is
port(
    
	CLK: in std_logic;
	D: in std_logic_vector(13 downto 0);
	RST: in std_logic;
	EN: in std_logic;
	Q: out std_logic_vector(13 downto 0)
	
	);
end ff_d_14;

architecture flipflop of ff_d_14 is
begin

	process(CLK, RST)
	begin
		if RST = '1' then
			Q <= "00000000000000";
		elsif (CLK'event and CLK = '1') then
			if EN = '1' then
				Q <= D;
			end if;
		end if;
	end process;	

end flipflop;